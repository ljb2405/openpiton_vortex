`include    "define.tmp.h"

`define NOC_DATA_BITS           `NOC_DATA_WIDTH-1:0