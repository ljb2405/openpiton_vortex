`include    "define.tmp.h"

`define NOC_DATA_BITS           `NOC_DATA_WIDTH-1:0
`define VORTEX_AXI_CTRL_ADDR_WIDTH  8
`define VORTEX_AXI_CTRL_DATA_WIDTH  32
`define VORTEX_AXI_MEM_ID_WIDTH 	32
`define VORTEX_AXI_MEM_ADDR_WIDTH   64
`define VORTEX_AXI_MEM_DATA_WIDTH   512