//`include  "define.tmp.h"

`define NOC_DATA_BITS                   `NOC_DATA_WIDTH-1:0
`define VX_DCR_ADDR_WIDTH               8
`define VX_DCR_DATA_WIDTH               32
`define VORTEX_AXI_MEM_ID_WIDTH 	    32
`define VORTEX_AXI_MEM_ADDR_WIDTH       64
`define VORTEX_AXI_MEM_DATA_WIDTH       512